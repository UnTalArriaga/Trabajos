LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ULTRASONICO IS
	PORT(
	CLK : IN STD_LOGIC;
	SENSOR_DISP : OUT STD_LOGIC;
	SENSOR_ECO : IN STD_LOGIC;
	SEGMENTOS : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
	SEGMENTOS2 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END ULTRASONICO;

ARCHITECTURE BEHAVIORAL OF ULTRASONICO IS
	FUNCTION NUMERO (DIGITO:UNSIGNED) RETURN STD_LOGIC_VECTOR IS
		VARIABLE HEX:STD_LOGIC_VECTOR(0 TO 7);
		BEGIN
			CASE DIGITO IS
				WHEN X"0" => HEX:="00000011";
				WHEN X"1" => HEX:="10011111";
				WHEN X"2" => HEX:="00100101";
				WHEN X"3" => HEX:="00001101";
				WHEN X"4" => HEX:="10011001";
				WHEN X"5" => HEX:="01001001";
				WHEN X"6" => HEX:="11000001";
				WHEN X"7" => HEX:="00011111";
				WHEN X"8" => HEX:="00000001";
				WHEN X"9" => HEX:="00001001";
				WHEN OTHERS => NULL;
			END CASE;
		RETURN(HEX);
	END NUMERO;
	
	SIGNAL CUENTA : UNSIGNED (16 DOWNTO 0) := (OTHERS => '0');
	SIGNAL CENTIMETROS : UNSIGNED (15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL CENTIMETROS_UNID : UNSIGNED (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL CENTIMETROS_DECE : UNSIGNED (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL SAL_UNID : UNSIGNED (3 DOWNTO 0) := (OTHERS => '0');	
	SIGNAL SAL_DECE : UNSIGNED (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL DIGITO : UNSIGNED (3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL ECO_PASADO : STD_LOGIC :='0';
	SIGNAL ECO_SINC : STD_LOGIC :='0';
	SIGNAL ECO_NSINC : STD_LOGIC :='0';
	SIGNAL ESPERA : STD_LOGIC :='0';
	SIGNAL SIETE_SEG_CUENTA : UNSIGNED (15 DOWNTO 0) := (OTHERS => '0');
	
BEGIN
	SIETE_SEG : PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF SIETE_SEG_CUENTA (SIETE_SEG_CUENTA'HIGH) = '1' THEN
				DIGITO <= SAL_UNID;
				SEGMENTOS <= NUMERO(DIGITO);
			ELSE
				DIGITO <= SAL_DECE;
				SEGMENTOS2 <= NUMERO(DIGITO);
			END IF;
			SIETE_SEG_CUENTA <= SIETE_SEG_CUENTA + 1;
		END IF;
		IF SAL_UNID < 10 AND SAL_DECE = 0 THEN
			SEGMENTOS2 <= "11111111";
			SEGMENTOS <= "01001001";
		END IF;
	END PROCESS;
	
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF ESPERA = '0' THEN
				IF CUENTA = 500 THEN
					SENSOR_DISP <= '0';
					ESPERA <= '1';
					CUENTA <= (OTHERS => '0');
				ELSE
					SENSOR_DISP <= '1';
					CUENTA <= CUENTA + 1;
				END IF;
			ELSIF ECO_PASADO = '0' AND ECO_SINC = '1' THEN
				CUENTA <= (OTHERS => '0');
				CENTIMETROS <= (OTHERS => '0');
				CENTIMETROS_UNID <= (OTHERS => '0');
				CENTIMETROS_DECE <= (OTHERS => '0');
			ELSIF ECO_PASADO = '1' AND ECO_SINC = '0' THEN
				SAL_UNID <= CENTIMETROS_UNID;
				SAL_DECE <= CENTIMETROS_DECE;
			ELSIF CUENTA = 2900-1 THEN
				IF CENTIMETROS_UNID = 9 THEN
					CENTIMETROS_UNID <= (OTHERS => '0');
					CENTIMETROS_DECE <= CENTIMETROS_DECE + 1;
				ELSE
					CENTIMETROS_UNID <= CENTIMETROS_UNID + 1;
				END IF;
				CENTIMETROS <= CENTIMETROS + 1;
				CUENTA <= (OTHERS => '0');
				IF CENTIMETROS = 3448 THEN
					ESPERA <= '0';
				END IF;
			ELSE
				CUENTA <= CUENTA + 1;
			END IF;
			ECO_PASADO <= ECO_SINC;
			ECO_SINC <= ECO_NSINC;
			ECO_NSINC <= SENSOR_ECO;
		END IF;
	END PROCESS;
END BEHAVIORAL;