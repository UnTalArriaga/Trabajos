LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MOTOR IS
	PORT(
		CLK : IN STD_LOGIC;
		DIR : IN STD_LOGIC;
		VEL : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		ACTIVO : IN STD_LOGIC;
		SALIDA : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END MOTOR;

ARCHITECTURE VELOCIDAD OF MOTOR IS
	SIGNAL STATE : STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL CONTADOR : INTEGER RANGE 0 TO 50000 := 0;
	SIGNAL TEMPORAL : STD_LOGIC;
	SIGNAL AUX1 : UNSIGNED (6 DOWNTO 0) := "1100100";
	SIGNAL CNT : UNSIGNED (6 DOWNTO 0);
	SIGNAL SALIDA_AUX : STD_LOGIC;
	
BEGIN
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF CONTADOR = 50000 THEN
				TEMPORAL <= NOT(TEMPORAL);
				CONTADOR <= 0;
			ELSE
				CONTADOR <= CONTADOR + 1;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (TEMPORAL, VEL)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF CNT = 99 THEN
				CNT <= (OTHERS => '0');
			ELSE
				CNT <= CNT + 1;
			END IF;
		END IF;
	END PROCESS;

	PROCESS (CLK)
	BEGIN
		IF VEL(0) = '1' THEN
			AUX1 <= "1100100";
		ELSIF VEL(1) = '1' THEN
			AUX1 <= "0110010";
		ELSIF VEL(2) = '1' THEN
			AUX1 <= "0001010";
		END IF;
	END PROCESS;
	
	SALIDA_AUX <= '1' WHEN (CNT < UNSIGNED (AUX1)) ELSE '0';
	
	PROCESS (TEMPORAL)
	BEGIN
		IF TEMPORAL'EVENT AND TEMPORAL = '1' THEN
			IF ACTIVO = '1' THEN
				IF DIR = '1' THEN
					STATE <= STATE + "01";
				END IF;
				IF DIR = '0' THEN
					STATE <= STATE - "01";
				END IF;
				CASE STATE IS
				WHEN "00" =>
					SALIDA(0) <= SALIDA_AUX;
					SALIDA(1) <= SALIDA_AUX;
					SALIDA(2) <= '0';
					SALIDA(3) <= '0';
				WHEN "01" =>
					SALIDA(0) <= '0';
					SALIDA(1) <= SALIDA_AUX;
					SALIDA(2) <= SALIDA_AUX;
					SALIDA(3) <= '0';
				WHEN "10" =>
					SALIDA(0) <= '0';
					SALIDA(1) <= '0';
					SALIDA(2) <= SALIDA_AUX;
					SALIDA(3) <= SALIDA_AUX;
				WHEN "11" =>
					SALIDA(0) <= SALIDA_AUX;
					SALIDA(1) <= '0';
					SALIDA(2) <= '0';
					SALIDA(3) <= SALIDA_AUX;
				END CASE;
			END IF;
		END IF;
	END PROCESS;
END VELOCIDAD;
	
	
	
	
	
	
	
	
	
	
	
	
	