LIBRARY IEEE;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LED IS
	PORT(
		CLK : IN STD_LOGIC;
		LED : OUT STD_LOGIC;
		ENTRADA : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		RESET : IN STD_LOGIC
	);
END LED;

ARCHITECTURE BEHAVIORAL OF LED IS
	SIGNAL CNT : UNSIGNED (6 DOWNTO 0);
BEGIN

	PROCESS (CLK, RESET, ENTRADA)
	BEGIN
		IF RESET = '1' THEN
			CNT <= (OTHERS => '0');
		ELSIF RISING_EDGE (CLK) THEN
			IF CNT = 99 THEN
				CNT <= (OTHERS => '0');
			ELSE
				CNT <= CNT + 1;
			END IF;
		END IF;
	END PROCESS;
	
	LED <= '1' WHEN (CNT < UNSIGNED(ENTRADA) ) ELSE '0';
END BEHAVIORAL;