LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY VGA IS
	GENERIC(
		CONSTANT H_PIXELS : INTEGER := 1024;
		CONSTANT H_FP : INTEGER := 8;
		CONSTANT H_PULSE : INTEGER := 176;
		CONSTANT H_BP : INTEGER := 56;
		
		CONSTANT V_PIXELS : INTEGER := 768;
		CONSTANT V_FP : INTEGER := 0;
		CONSTANT V_PULSE : INTEGER := 8;
		CONSTANT V_BP : INTEGER := 41
	);
	PORT(
		CLK : IN STD_LOGIC;
		RED : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		GREEN : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		BLUE : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		H_SYNC : OUT STD_LOGIC;
		V_SYNC : OUT STD_LOGIC
	);
END VGA;

ARCHITECTURE BEHAVIORAL OF VGA IS
	SIGNAL H_PERIOD : INTEGER := H_PULSE + H_BP + H_PIXELS + H_FP;
	SIGNAL V_PERIOD : INTEGER := V_PULSE + V_BP + V_PIXELS + V_FP;
	SIGNAL H_COUNT : INTEGER RANGE 0 TO H_PERIOD - 1 := 0;
	SIGNAL V_COUNT : INTEGER RANGE 0 TO V_PERIOD - 1 := 0;
	SIGNAL RELOJ_PIXEL : STD_LOGIC;
	SIGNAL COLUMN : INTEGER RANGE 0 TO H_PERIOD - 1 := 0;
	SIGNAL ROW : INTEGER RANGE 0 TO V_PERIOD - 1 := 0;
	SIGNAL DISPLAY_ENA : STD_LOGIC;
	
BEGIN
	PROCESS (CLK)
	BEGIN
		RELOJ_PIXEL <= CLK;
	END PROCESS;
	
	PROCESS (RELOJ_PIXEL)
	BEGIN
		IF RISING_EDGE(RELOJ_PIXEL) THEN
			IF H_COUNT < H_PERIOD - 1 THEN
				H_COUNT <= H_COUNT + 1;
			ELSE
				H_COUNT <= 0;
				IF V_COUNT < V_PERIOD - 1 THEN
					V_COUNT <= V_COUNT + 1;
				ELSE
					V_COUNT <= 0;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (RELOJ_PIXEL)
	BEGIN
		IF RISING_EDGE(RELOJ_PIXEL) THEN
			IF H_COUNT > (H_PIXELS + H_FP) OR H_COUNT > (H_PIXELS + H_FP + H_PULSE) THEN
				H_SYNC <= '0';
			ELSE
				H_SYNC <= '1';
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (RELOJ_PIXEL)
	BEGIN
		IF RISING_EDGE(RELOJ_PIXEL) THEN
			IF V_COUNT > (V_PIXELS + V_FP) OR V_COUNT > (V_PIXELS + V_FP + V_PULSE) THEN
				V_SYNC <= '0';
			ELSE
				V_SYNC <= '1';
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (RELOJ_PIXEL)
	BEGIN
		IF RISING_EDGE(RELOJ_PIXEL) THEN
			IF H_COUNT < H_PIXELS THEN
				COLUMN <= H_COUNT;
			END IF;
			IF V_COUNT < V_PIXELS THEN
				ROW <= V_COUNT;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (RELOJ_PIXEL)
	BEGIN
		IF RISING_EDGE(RELOJ_PIXEL) THEN
			IF H_COUNT < H_PIXELS AND V_COUNT < V_PIXELS THEN
				DISPLAY_ENA <= '1';
			ELSE
				DISPLAY_ENA <= '0';
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS (DISPLAY_ENA, ROW, COLUMN)
	BEGIN
		IF DISPLAY_ENA = '1' THEN
			IF ((ROW > 300 AND ROW < 350) AND (COLUMN > 350 AND COLUMN < 400)) THEN
				RED <= (OTHERS => '1');
				GREEN <= (OTHERS => '1');
				BLUE <= (OTHERS => '0');
			ELSIF ((ROW > 300 AND ROW < 350) AND (COLUMN > 450 AND COLUMN < 500)) THEN
				RED <= (OTHERS => '0');
				GREEN <= (OTHERS => '1');
				BLUE <= (OTHERS => '1');
			ELSIF ((ROW > 300 AND ROW < 350) AND (COLUMN > 550 AND COLUMN < 600)) THEN
				RED <= (OTHERS => '1');
				GREEN <= (OTHERS => '1');
				BLUE <= (OTHERS => '1');
			END IF;
		ELSE
			RED <= (OTHERS => '0');
			GREEN <= (OTHERS => '0');
			BLUE <= (OTHERS => '0');
		END IF;
	END PROCESS;
END BEHAVIORAL;
	
	
	